module nandg(output Y, input A, B);
    nand(Y, A, B); 
endmodule
