// Code your design here
module org(output Y, input A, B);
    or(Y, A, B); 
endmodule
