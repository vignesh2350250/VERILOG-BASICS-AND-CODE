// Code your design here
module andg(output A, input B, Y);
  and(A, B, Y); 
endmodule
