module xorg(input A, B, output Y);
  xor(Y,A,B);
endmodule 

  
