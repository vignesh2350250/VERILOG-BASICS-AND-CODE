class transaction;
  bit clk;
  bit rst;
  bit [8:0]addr;
  bit [8:0]data;
  bit we;
  bit re;
  reg [8:0]datao;
  
endclass
  
  
