interface operation;
  logic clk,rst,d;
  logic q;
endinterface
