class transaction;
  bit clk;
  bit rst;
 reg d;
  bit q;
endclass
  
  
