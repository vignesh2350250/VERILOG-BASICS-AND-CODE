interface operation;
  logic clk,rst;
  logic [8:0]data;
  logic [8:0]addr;
  logic we,re;
  logic [8:0]datao;
endinterface
