class transaction;
  bit clk;
  rand bit rst;
  bit en;
  bit ds;
  reg [7:0]ctr;
endclass
