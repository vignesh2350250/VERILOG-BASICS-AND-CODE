module norg(input A, B ,output Y);
  nor(Y,A,B);
endmodule
  
