interface inter;
  logic clk;
  logic rst;
  logic en;
  logic ds;
  logic [7:0]ctr;
endinterface
