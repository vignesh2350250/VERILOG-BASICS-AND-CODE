module andg(output z, input x, y);
  and(z, x, y); 
endmodule
